library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Mini_projecto_fase3 is
	port(SW                             : in std_logic_vector(1 downto 0);
		  CLOCK_50                       : in std_logic;
		  KEY                            : in std_logic_vector(3 downto 0);
		  HEX0, HEX1,HEX2,HEX3,HEX4,HEX5 : out std_logic_vector(6 downto 0);
		  LEDG                           : out std_logic_vector(8 downto 0));
end Mini_projecto_fase3;

architecture SHell of Mini_projecto_fase3 is

	signal s_clk1Hz, s_clk4Hz, s_termCount, s_hex0En, s_hex1En, s_hex5En, s_hex4En, s_hex3En, s_setM, s_setS, s_set : std_logic;
	signal s_hex2, s_hex3, s_hex4, s_hex5 : std_logic_vector(4 downto 0);
	signal s_count  : std_logic_vector(15 downto 0);

begin

	clk1Hz  : entity work.ClkDividerN(RTL)
						generic map(k => 50000000)
						port map(clkIn  => CLOCK_50,
									clkOut => s_clk1Hz);
					
	clk4Hz  : entity work.ClkDividerN(RTL)
						generic map(k => 12500000)
						port map(clkIn  => CLOCK_50,
									clkOut => s_clk4Hz);
									
	s_setM <= (not KEY(2)) and (not KEY(3));	
	s_setS <= (not KEY(2)) and (not KEY(1));	
	s_set  <= not KEY(2);								
	
	Counter : entity work.TimerCounter(Behavioral)
						port map(clk       => s_clk1Hz,
									clkSet    => s_clk4Hz,
									set       => s_set,
									setM      => s_setM,
									setS      => s_setS,
									enable    => SW(0),
									reset     => SW(1),
									start     => key(0),
									countOut  => s_count,
									termCount => s_termCount);
									
	s_hex2 <= ('0' & s_count(3 downto 0)) when (s_termCount = '0') else "00001";
	s_hex3 <= ('0' & s_count(7 downto 4)) when (s_termCount = '0') else "10001";
	s_hex4 <= ('0' & s_count(11 downto 8)) when (s_termCount = '0') else "00001";
	s_hex5 <= ('0' & s_count(15 downto 12)) when (s_termCount = '0') else "01111";
	
	s_hex0En <= s_termCount;
	s_hex1En <= s_termCount;
	s_hex5En <= '1' when (s_count(15 downto 12) /= x"0" or s_termCount = '1') else '0';
	s_hex4En <= '1' when (s_count(15 downto 8) /= x"00" or s_termCount = '1') else '0';
	s_hex3En <= '1' when (s_count(15 downto 4) /= x"000" or s_termCount = '1') else '0';
							
	Hex0Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => "10010",
									enable   => s_hex0En,
									decOut_n => HEX0);
			
	Hex1Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => "00101",
									enable   => s_hex1En,
									decOut_n => HEX1);
									
	Hex2Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => s_hex2,
									enable   => '1',
									decOut_n => HEX2);								
	
	
	Hex3Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => s_hex3,
									enable   => s_hex3En,
									decOut_n => HEX3);
	
	Hex4Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => s_hex4,
									enable   => s_hex4En,
									decOut_n => HEX4);	
									
	Hex5Dec    : entity work.Bin7SegDecoder(Behavioral)
						port map(binInput => s_hex5,
									enable   => s_hex5En,
									decOut_n => HEX5);
			
	LEDG(8) <= s_clk1Hz and (not s_termCount);
	
end Shell;